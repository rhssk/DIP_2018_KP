-- library IEEE;
-- use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

-- entity TOP0 is
-- end TOP0;

-- architecture Behavioral of TOP0 is

-- begin


-- end Behavioral;
